module set_clock1 (output reg [3:0] s1h0 = 0, s1h1 = 0, s1m0 = 0, s1m1 = 0,
						input switch,
						input reset,
						input push2, push3
						);	

// Set minute						
always @(posedge reset, negedge push2) begin
	if (reset == 1) begin
			s1m0 <= 0;
			s1m1 <= 0;
	end
	else begin
		if ( (push2 == 0) ) begin
			if(switch == 1) begin
				if ((s1m0 < 4'd9)) begin
					s1m0 <= s1m0 + 1;
					s1m1 <= s1m1;
				end
				else begin
					s1m0 <= 0;
					if (s1m1 < 4'd5)
						s1m1 <= s1m1 + 1;
					else 
						s1m1 <= 0;
				end
			end
			else begin
				s1m0<= s1m0;
				s1m1<= s1m1;
			end
		end
		else begin
	
			s1m0 <= s1m0;
			s1m1 <= s1m1;

		end
	end
end

// Set hour
always@(posedge reset, negedge push3) begin
	if (reset == 1) begin
		s1h0 <= 0;
		s1h1 <= 0; 
	end
	else begin
		if(push3 == 0) begin
			if(switch == 1) begin
				if ( (s1h1 <= 4'd1) && ( s1h0 < 4'd9) )
					s1h0 <= s1h0 + 1;
				else if ( (s1h1 == 4'd2) && ( s1h0 < 4'd3) )
					s1h0 <= s1h0 + 1;
				else begin
					s1h0 <= 0;
					if (s1h1 < 4'd2)
						s1h1 <= s1h1 + 1;
					else 
						s1h1 <= 4'd0;
				end
			end
			else begin
				s1h0 <= s1h0;
				s1h1 <= s1h1;
			end
		end 
		else begin
			s1h0 <= s1h0;
			s1h1 <= s1h1; 
		end 	
	end 
end 
	
endmodule
